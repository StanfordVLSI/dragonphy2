module input_buffer (
	input inp,
	input inm,
	input pd,
	output clk
);
endmodule
