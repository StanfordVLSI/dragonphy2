module MOMcap (
    input Ctop,
    output Cbot
);
endmodule


