`ifndef INIT_EXT_PI_CODE
	`define INIT_EXT_PI_CODE 'd0
`endif

`default_nettype none

module adbg_stim import const_pack::*; (
	acore_debug_intf adbg_intf_i
);




endmodule

`default_nettype wire