
module inv_3_fixed (input in, output out );
assign out = ~(in);
endmodule

