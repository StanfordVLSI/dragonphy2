
module inv_v2t_5_fixed (input in, output out );
assign out = ~(in);
endmodule

