module CS_cell_dmm ();
endmodule


