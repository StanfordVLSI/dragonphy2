module ff_c_sn_rn(
    input D,
    input CP,
    input CDN,
    output Q
);
endmodule
