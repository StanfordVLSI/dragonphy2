module vio (
    output wire logic emu_rst,
    input wire logic [63:0] number,
    input wire logic clk
);

    // instantiate vio here...

endmodule
