`ifndef __VOLTAGE_NET_SV__
`define __VOLTAGE_NET_SV__
`endif // `ifndef __VOLTAGE_NET_SV__
