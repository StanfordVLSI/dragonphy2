
module SW (input IN, input CLK, input CLKB, output OUT);
endmodule


