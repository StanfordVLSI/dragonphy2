* Automatically generated file.
.include /home/dstanley/research/dragonphy/model_generation/comparator/comparator.sp
X0 my_in my_out vdd vss simple_comparator
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    Gs sw_p sw_n cur='V(sw_p, sw_n)*(0.999999999*V(ctl_p, ctl_n)+1e-09)'
.ends
X1 __vdd_v vdd __vdd_s 0 inout_sw_mod
V2 __vdd_v 0 DC 1.2 PWL(0 1.2 2.6000000000000016e-07 1.2)
V3 __vdd_s 0 DC 1 PWL(0 1 2.6000000000000016e-07 1)
X4 __vss_v vss __vss_s 0 inout_sw_mod
V5 __vss_v 0 DC 0 PWL(0 0 5e-09 0 5.2e-09 0.0 2.6000000000000016e-07 0.0)
V6 __vss_s 0 DC 1 PWL(0 1 5e-09 1 5.2e-09 1 2.6000000000000016e-07 1)
X7 __my_in_v my_in __my_in_s 0 inout_sw_mod
V8 __my_in_v 0 DC 0 PWL(0 0 1e-08 0 1.02e-08 0.0013793424693735947 1.5000000000000002e-08 0.0013793424693735947 1.52e-08 0.025846956206025992 2e-08 0.025846956206025992 2.02e-08 0.055839779183417176 2.5e-08 0.055839779183417176 2.5199999999999997e-08 0.08019992204882016 3e-08 0.08019992204882016 3.02e-08 0.11070028793547686 3.4999999999999996e-08 0.11070028793547686 3.52e-08 0.12371380601275465 3.9999999999999994e-08 0.12371380601275465 4.0199999999999996e-08 0.1473347937622795 4.499999999999999e-08 0.1473347937622795 4.5199999999999994e-08 0.17909547788612704 4.999999999999999e-08 0.17909547788612704 5.019999999999999e-08 0.20267662263598074 5.499999999999999e-08 0.20267662263598074 5.519999999999999e-08 0.2356081371884854 6e-08 0.2356081371884854 6.02e-08 0.244463774582808 6.5e-08 0.244463774582808 6.52e-08 0.28340259247220917 7e-08 0.28340259247220917 7.02e-08 0.29198563988220183 7.500000000000001e-08 0.29198563988220183 7.520000000000001e-08 0.3125544775385783 8.000000000000001e-08 0.3125544775385783 8.020000000000002e-08 0.34468981539054766 8.500000000000002e-08 0.34468981539054766 8.520000000000002e-08 0.37199395148667186 9.000000000000003e-08 0.37199395148667186 9.020000000000003e-08 0.4038357186906867 9.500000000000003e-08 0.4038357186906867 9.520000000000003e-08 0.41471533451865045 1.0000000000000004e-07 0.41471533451865045 1.0020000000000004e-07 0.4410140366180115 1.0500000000000004e-07 0.4410140366180115 1.0520000000000004e-07 0.4674401669937914 1.1000000000000005e-07 0.4674401669937914 1.1020000000000005e-07 0.49778503095477666 1.1500000000000005e-07 0.49778503095477666 1.1520000000000005e-07 0.5104127487210219 1.2000000000000004e-07 0.5104127487210219 1.2020000000000003e-07 0.5504008080749023 1.2500000000000005e-07 0.5504008080749023 1.2520000000000004e-07 0.562279014136317 1.3000000000000005e-07 0.562279014136317 1.3020000000000004e-07 0.5857031766911577 1.3500000000000006e-07 0.5857031766911577 1.3520000000000005e-07 0.6204235103891967 1.4000000000000006e-07 0.6204235103891967 1.4020000000000005e-07 0.6333717934759027 1.4500000000000007e-07 0.6333717934759027 1.4520000000000006e-07 0.6533594260369466 1.5000000000000007e-07 0.6533594260369466 1.5020000000000006e-07 0.6872138380598609 1.5500000000000008e-07 0.6872138380598609 1.5520000000000007e-07 0.7000106084426347 1.6000000000000008e-07 0.7000106084426347 1.6020000000000007e-07 0.7207562016367184 1.650000000000001e-07 0.7207562016367184 1.6520000000000008e-07 0.7468160898459608 1.700000000000001e-07 0.7468160898459608 1.7020000000000008e-07 0.7851958420721956 1.750000000000001e-07 0.7851958420721956 1.7520000000000009e-07 0.8045253018773233 1.800000000000001e-07 0.8045253018773233 1.802000000000001e-07 0.8307772158277528 1.850000000000001e-07 0.8307772158277528 1.852000000000001e-07 0.8427691909806514 1.900000000000001e-07 0.8427691909806514 1.902000000000001e-07 0.8678196828992881 1.9500000000000012e-07 0.8678196828992881 1.952000000000001e-07 0.9048672615938991 2.0000000000000012e-07 0.9048672615938991 2.002000000000001e-07 0.9221454803476127 2.0500000000000013e-07 0.9221454803476127 2.0520000000000012e-07 0.9388985083012233 2.1000000000000013e-07 0.9388985083012233 2.1020000000000012e-07 0.9720012036386739 2.1500000000000014e-07 0.9720012036386739 2.1520000000000013e-07 0.9993916986343694 2.2000000000000014e-07 0.9993916986343694 2.2020000000000013e-07 1.0091848616677421 2.2500000000000015e-07 1.0091848616677421 2.2520000000000014e-07 1.0471412012594195 2.3000000000000015e-07 1.0471412012594195 2.3020000000000014e-07 1.068035524340207 2.3500000000000016e-07 1.068035524340207 2.3520000000000015e-07 1.0823645072107246 2.4000000000000014e-07 1.0823645072107246 2.4020000000000015e-07 1.105981285973563 2.4500000000000014e-07 1.105981285973563 2.4520000000000016e-07 1.1337153045653219 2.5000000000000015e-07 1.1337153045653219 2.5020000000000016e-07 1.1561545467385101 2.5500000000000015e-07 1.1561545467385101 2.5520000000000017e-07 1.1780933382308891 2.6000000000000016e-07 1.1780933382308891)
V9 __my_in_s 0 DC 1 PWL(0 1 1e-08 1 1.02e-08 1 1.5000000000000002e-08 1 1.52e-08 1 2e-08 1 2.02e-08 1 2.5e-08 1 2.5199999999999997e-08 1 3e-08 1 3.02e-08 1 3.4999999999999996e-08 1 3.52e-08 1 3.9999999999999994e-08 1 4.0199999999999996e-08 1 4.499999999999999e-08 1 4.5199999999999994e-08 1 4.999999999999999e-08 1 5.019999999999999e-08 1 5.499999999999999e-08 1 5.519999999999999e-08 1 6e-08 1 6.02e-08 1 6.5e-08 1 6.52e-08 1 7e-08 1 7.02e-08 1 7.500000000000001e-08 1 7.520000000000001e-08 1 8.000000000000001e-08 1 8.020000000000002e-08 1 8.500000000000002e-08 1 8.520000000000002e-08 1 9.000000000000003e-08 1 9.020000000000003e-08 1 9.500000000000003e-08 1 9.520000000000003e-08 1 1.0000000000000004e-07 1 1.0020000000000004e-07 1 1.0500000000000004e-07 1 1.0520000000000004e-07 1 1.1000000000000005e-07 1 1.1020000000000005e-07 1 1.1500000000000005e-07 1 1.1520000000000005e-07 1 1.2000000000000004e-07 1 1.2020000000000003e-07 1 1.2500000000000005e-07 1 1.2520000000000004e-07 1 1.3000000000000005e-07 1 1.3020000000000004e-07 1 1.3500000000000006e-07 1 1.3520000000000005e-07 1 1.4000000000000006e-07 1 1.4020000000000005e-07 1 1.4500000000000007e-07 1 1.4520000000000006e-07 1 1.5000000000000007e-07 1 1.5020000000000006e-07 1 1.5500000000000008e-07 1 1.5520000000000007e-07 1 1.6000000000000008e-07 1 1.6020000000000007e-07 1 1.650000000000001e-07 1 1.6520000000000008e-07 1 1.700000000000001e-07 1 1.7020000000000008e-07 1 1.750000000000001e-07 1 1.7520000000000009e-07 1 1.800000000000001e-07 1 1.802000000000001e-07 1 1.850000000000001e-07 1 1.852000000000001e-07 1 1.900000000000001e-07 1 1.902000000000001e-07 1 1.9500000000000012e-07 1 1.952000000000001e-07 1 2.0000000000000012e-07 1 2.002000000000001e-07 1 2.0500000000000013e-07 1 2.0520000000000012e-07 1 2.1000000000000013e-07 1 2.1020000000000012e-07 1 2.1500000000000014e-07 1 2.1520000000000013e-07 1 2.2000000000000014e-07 1 2.2020000000000013e-07 1 2.2500000000000015e-07 1 2.2520000000000014e-07 1 2.3000000000000015e-07 1 2.3020000000000014e-07 1 2.3500000000000016e-07 1 2.3520000000000015e-07 1 2.4000000000000014e-07 1 2.4020000000000015e-07 1 2.4500000000000014e-07 1 2.4520000000000016e-07 1 2.5000000000000015e-07 1 2.5020000000000016e-07 1 2.5500000000000015e-07 1 2.5520000000000017e-07 1 2.6000000000000016e-07 1)
.probe my_out
.ic
.tran 2.6000000000000014e-10 2.6000000000000016e-07
.control
run
set filetype=ascii
write
exit
.endc
.end
