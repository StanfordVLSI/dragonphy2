
module inv_v2t_2_fixed (input in, output out );
assign out = ~(in);
endmodule

