`ifndef __IOTYPE_SV__
`define __IOTYPE_SV__

    `include "mLingua_pwl.vh"
    `include "voltage_net.sv"
    
    `define pwl_t pwl
    `define real_t real
    `define voltage_t wire
    
    `define PWL_ZERO '{0,0,0}

`endif // `ifndef __IOTYPE_SV__
