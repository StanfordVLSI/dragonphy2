module inv_2 (
    input in,
    output out
);
endmodule

