
module inv_gf (input in, output out );
assign out = ~(in);
endmodule

