module input_buffer (
	input inp,
	input inm,
	input pd,
	output clk,
	output clk_b
);
endmodule
