
module inv_bld_4_fixed (input in, output out );
assign out = ~(in);
endmodule

