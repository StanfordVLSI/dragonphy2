`ifndef __IOTYPE_SV__
`define __IOTYPE_SV__

    `include "mLingua_pwl.vh"

    `define pwl_t pwl
    `define real_t real
    `define voltage_t real

    `define PWL_ZERO '{0,0,0}
    `define SIMULATION

`endif // `ifndef __IOTYPE_SV__
