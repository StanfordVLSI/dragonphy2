`ifndef __IOTYPE_SV__
`define __IOTYPE_SV__

    `define pwl_t wire logic [15:0]
	`define real_t wire logic
	`define voltage_t wire logic

	`define PWL_ZERO 1'b0

`endif // `ifndef __IOTYPE_SV__
