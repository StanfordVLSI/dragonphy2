/********************************************************************
filename: phase_blender.sv

Description: 
multi-bit phase blender.

Assumptions:

Todo:

********************************************************************/

`include "mLingua_pwl.vh"

`default_nettype none

module phase_blender import const_pack::*; #(
// parameters here
  parameter integer Nblender = 4,  // # of control bit
  parameter real del_nom = 100e-12, // intrinsic delay
  parameter real del_std = 0e-12,
  parameter real jit_rms = 0e-15
) (
// I/Os here
    input wire logic [1:0]  ph_in,                  // two clocks being interpolated
    input wire logic [2**Nblender-1:0] sel_bld_thm, // interpolation weight (thermometer coded) 
    output reg ph_out                               // blended clock
);

timeunit 1fs;
timeprecision 1fs;

real TU = 1/1s; // verilog time unit in sec

//----- VARIABLE/SIGNAL DECLARATION -----
integer sel_bld_bin;    // binary value of sel_bld_thm
real t_lead;
real tdiff; // time difference b/t two clock phases
real tout;  // phase interpolated delay
real wgt;       // phase interpolation weight
real td, rj;    // delay of this cell, random jitter
logic sign;     // indicates which clock leads the other
logic ph_lead;  // selected clock that leads the other
logic ph_in0_d, ph_in1_d;   // delayed signal of ph_in[0], ph_in[1]
real lut [17];  // interpolation weight LUT

initial begin
    lut[0]=0.0;
    lut[1]=0.0625;
    lut[2]=0.125;
    lut[3]=0.1875;
    lut[4]=0.25;
    lut[5]=0.3125;
    lut[6]=0.375;
    lut[7]=0.4375;
    lut[8]=0.5;
    lut[9]=0.5625;
    lut[10]=0.625;
    lut[11]=0.6875;
    lut[12]=0.75;
    lut[13]=0.8125;
    lut[14]=0.875;
    lut[15]=0.9375;
    lut[16]=1.0;
end


//----- FUNCTIONAL DESCRIPTION -----

// design parameter class init
PIParameter pi_obj;

initial begin
    pi_obj = new();
    td = pi_obj.td_mixermb;
end

// phase interpolation weight
assign sel_bld_bin = $countones(sel_bld_thm) ;

`ifdef LUT
    assign wgt = real'(lut[sel_bld_bin]) ;
`else
    assign wgt = real'(sel_bld_bin)/2.0**Nblender ;
`endif

// delay two inputs
always @(ph_in[0])  ph_in0_d <= #(td*1s) ph_in[0];
always @(ph_in[1])  ph_in1_d <= #(td*1s) ph_in[1];

// find which clock input leads
always @(ph_in[0])  sign <= ph_in[0] ^ ph_in[1];
assign ph_lead = sign ? ph_in0_d : ph_in1_d; 

// compute the phase difference
always @(ph_in) begin
    if (ph_in[0] ^ ph_in[1]) 
        t_lead = `get_time;
    else begin
        tdiff = `get_time - t_lead;
        tout = tdiff * wgt;
    end
end

// phase interpolation
always @(*) begin
    rj = pi_obj.get_rj_mixermb();
    if (sign)   ph_out <= `delay(tout+rj)       ph_in0_d;
    else        ph_out <= `delay(tdiff-tout+rj) ph_in1_d;
end


//always @(del, td, jit) begin
//	assert ( Nblender==0 || del+jit > td || $realtime*TU < 100e-9 ) else $warning("%m: del+jit (%f [psec]) is less than td(%f [psec]) at %f [nsec]", (del+jit)/1e-12, td/1e-12, $realtime*TU*1e9);
//end

endmodule

`default_nettype wire
