package constant_pack;
	localparam integer channel_width = 16;
	localparam integer code_precision = 8;
	localparam integer ffe_length = 5;
	localparam integer ffe_weight_precision = 8;
endpackage
