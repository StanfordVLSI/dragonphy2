* Automatically generated file.
.include /home/dstanley/research/dragonphy/model_generation/comparator.sp
X0 my_in my_out vdd vss simple_comparator
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    Gs sw_p sw_n cur='V(sw_p, sw_n)*(0.999999999*V(ctl_p, ctl_n)+1e-09)'
.ends
X1 __vdd_v vdd __vdd_s 0 inout_sw_mod
V2 __vdd_v 0 DC 1.2 PWL(0 1.2 2.6000000000000016e-07 1.2)
V3 __vdd_s 0 DC 1 PWL(0 1 2.6000000000000016e-07 1)
X4 __vss_v vss __vss_s 0 inout_sw_mod
V5 __vss_v 0 DC 0 PWL(0 0 5e-09 0 5.2e-09 0.0 2.6000000000000016e-07 0.0)
V6 __vss_s 0 DC 1 PWL(0 1 5e-09 1 5.2e-09 1 2.6000000000000016e-07 1)
X7 __my_in_v my_in __my_in_s 0 inout_sw_mod
V8 __my_in_v 0 DC 0 PWL(0 0 1e-08 0 1.02e-08 0.01545130023088627 1.5000000000000002e-08 0.01545130023088627 1.52e-08 0.02898629045640844 2e-08 0.02898629045640844 2.02e-08 0.052663059550690165 2.5e-08 0.052663059550690165 2.5199999999999997e-08 0.09108106205162704 3e-08 0.09108106205162704 3.02e-08 0.11388070818919939 3.4999999999999996e-08 0.11388070818919939 3.52e-08 0.1333307057693876 3.9999999999999994e-08 0.1333307057693876 4.0199999999999996e-08 0.15454110931443513 4.499999999999999e-08 0.15454110931443513 4.5199999999999994e-08 0.1807224256043586 4.999999999999999e-08 0.1807224256043586 5.019999999999999e-08 0.1934821071385532 5.499999999999999e-08 0.1934821071385532 5.519999999999999e-08 0.2347108595955626 6e-08 0.2347108595955626 6.02e-08 0.24387954619221064 6.5e-08 0.24387954619221064 6.52e-08 0.2720283371965442 7e-08 0.2720283371965442 7.02e-08 0.30425614474474594 7.500000000000001e-08 0.30425614474474594 7.520000000000001e-08 0.3299213446264103 8.000000000000001e-08 0.3299213446264103 8.020000000000002e-08 0.3527607374124997 8.500000000000002e-08 0.3527607374124997 8.520000000000002e-08 0.3606022205821702 9.000000000000003e-08 0.3606022205821702 9.020000000000003e-08 0.38986714447869125 9.500000000000003e-08 0.38986714447869125 9.520000000000003e-08 0.4293423036336924 1.0000000000000004e-07 0.4293423036336924 1.0020000000000004e-07 0.45392883985042753 1.0500000000000004e-07 0.45392883985042753 1.0520000000000004e-07 0.4686047241506314 1.1000000000000005e-07 0.4686047241506314 1.1020000000000005e-07 0.49585802632395864 1.1500000000000005e-07 0.49585802632395864 1.1520000000000005e-07 0.5125469564735915 1.2000000000000004e-07 0.5125469564735915 1.2020000000000003e-07 0.5344720082726491 1.2500000000000005e-07 0.5344720082726491 1.2520000000000004e-07 0.5656088673564488 1.3000000000000005e-07 0.5656088673564488 1.3020000000000004e-07 0.5838735582271181 1.3500000000000006e-07 0.5838735582271181 1.3520000000000005e-07 0.6195621745725977 1.4000000000000006e-07 0.6195621745725977 1.4020000000000005e-07 0.6438945945105092 1.4500000000000007e-07 0.6438945945105092 1.4520000000000006e-07 0.659903310004599 1.5000000000000007e-07 0.659903310004599 1.5020000000000006e-07 0.6735460116950088 1.5500000000000008e-07 0.6735460116950088 1.5520000000000007e-07 0.7150735699119537 1.6000000000000008e-07 0.7150735699119537 1.6020000000000007e-07 0.7301361952618605 1.650000000000001e-07 0.7301361952618605 1.6520000000000008e-07 0.7628747971316017 1.700000000000001e-07 0.7628747971316017 1.7020000000000008e-07 0.7693369310696362 1.750000000000001e-07 0.7693369310696362 1.7520000000000009e-07 0.802786541738852 1.800000000000001e-07 0.802786541738852 1.802000000000001e-07 0.8280532706974941 1.850000000000001e-07 0.8280532706974941 1.852000000000001e-07 0.8480662974745661 1.900000000000001e-07 0.8480662974745661 1.902000000000001e-07 0.8651422620766508 1.9500000000000012e-07 0.8651422620766508 1.952000000000001e-07 0.9106671271560167 2.0000000000000012e-07 0.9106671271560167 2.002000000000001e-07 0.9342854042604054 2.0500000000000013e-07 0.9342854042604054 2.0520000000000012e-07 0.9360165891041062 2.1000000000000013e-07 0.9360165891041062 2.1020000000000012e-07 0.9632616019095865 2.1500000000000014e-07 0.9632616019095865 2.1520000000000013e-07 1.0055782396500856 2.2000000000000014e-07 1.0055782396500856 2.2020000000000013e-07 1.011784036251235 2.2500000000000015e-07 1.011784036251235 2.2520000000000014e-07 1.0526114984511517 2.3000000000000015e-07 1.0526114984511517 2.3020000000000014e-07 1.0562507068869527 2.3500000000000016e-07 1.0562507068869527 2.3520000000000015e-07 1.088300167949501 2.4000000000000014e-07 1.088300167949501 2.4020000000000015e-07 1.1239462360933608 2.4500000000000014e-07 1.1239462360933608 2.4520000000000016e-07 1.146116105030656 2.5000000000000015e-07 1.146116105030656 2.5020000000000016e-07 1.1547314347180633 2.5500000000000015e-07 1.1547314347180633 2.5520000000000017e-07 1.1957696805729963 2.6000000000000016e-07 1.1957696805729963)
V9 __my_in_s 0 DC 1 PWL(0 1 1e-08 1 1.02e-08 1 1.5000000000000002e-08 1 1.52e-08 1 2e-08 1 2.02e-08 1 2.5e-08 1 2.5199999999999997e-08 1 3e-08 1 3.02e-08 1 3.4999999999999996e-08 1 3.52e-08 1 3.9999999999999994e-08 1 4.0199999999999996e-08 1 4.499999999999999e-08 1 4.5199999999999994e-08 1 4.999999999999999e-08 1 5.019999999999999e-08 1 5.499999999999999e-08 1 5.519999999999999e-08 1 6e-08 1 6.02e-08 1 6.5e-08 1 6.52e-08 1 7e-08 1 7.02e-08 1 7.500000000000001e-08 1 7.520000000000001e-08 1 8.000000000000001e-08 1 8.020000000000002e-08 1 8.500000000000002e-08 1 8.520000000000002e-08 1 9.000000000000003e-08 1 9.020000000000003e-08 1 9.500000000000003e-08 1 9.520000000000003e-08 1 1.0000000000000004e-07 1 1.0020000000000004e-07 1 1.0500000000000004e-07 1 1.0520000000000004e-07 1 1.1000000000000005e-07 1 1.1020000000000005e-07 1 1.1500000000000005e-07 1 1.1520000000000005e-07 1 1.2000000000000004e-07 1 1.2020000000000003e-07 1 1.2500000000000005e-07 1 1.2520000000000004e-07 1 1.3000000000000005e-07 1 1.3020000000000004e-07 1 1.3500000000000006e-07 1 1.3520000000000005e-07 1 1.4000000000000006e-07 1 1.4020000000000005e-07 1 1.4500000000000007e-07 1 1.4520000000000006e-07 1 1.5000000000000007e-07 1 1.5020000000000006e-07 1 1.5500000000000008e-07 1 1.5520000000000007e-07 1 1.6000000000000008e-07 1 1.6020000000000007e-07 1 1.650000000000001e-07 1 1.6520000000000008e-07 1 1.700000000000001e-07 1 1.7020000000000008e-07 1 1.750000000000001e-07 1 1.7520000000000009e-07 1 1.800000000000001e-07 1 1.802000000000001e-07 1 1.850000000000001e-07 1 1.852000000000001e-07 1 1.900000000000001e-07 1 1.902000000000001e-07 1 1.9500000000000012e-07 1 1.952000000000001e-07 1 2.0000000000000012e-07 1 2.002000000000001e-07 1 2.0500000000000013e-07 1 2.0520000000000012e-07 1 2.1000000000000013e-07 1 2.1020000000000012e-07 1 2.1500000000000014e-07 1 2.1520000000000013e-07 1 2.2000000000000014e-07 1 2.2020000000000013e-07 1 2.2500000000000015e-07 1 2.2520000000000014e-07 1 2.3000000000000015e-07 1 2.3020000000000014e-07 1 2.3500000000000016e-07 1 2.3520000000000015e-07 1 2.4000000000000014e-07 1 2.4020000000000015e-07 1 2.4500000000000014e-07 1 2.4520000000000016e-07 1 2.5000000000000015e-07 1 2.5020000000000016e-07 1 2.5500000000000015e-07 1 2.5520000000000017e-07 1 2.6000000000000016e-07 1)
.probe my_out
.ic
.tran 2.6000000000000014e-10 2.6000000000000016e-07
.control
run
set filetype=ascii
write
exit
.endc
.end
