module biasgen import const_pack::Nbias; (
    input en,
    input [Nbias-1:0] ctl,
    input Vbias
);
endmodule
