module tri_buff_fixed (
    input in,
    input en,
    output out
);

bufif1(out,in,en);

endmodule




