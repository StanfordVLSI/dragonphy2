`ifndef __SIGNALS_SV__
`define __SIGNALS_SV__

`define ANALOG_INPUT inout wire
`define ANALOG_OUTPUT inout wire

`define DECL_ANALOG(x) wire x;

`endif // `ifndef __SIGNALS_SV__
