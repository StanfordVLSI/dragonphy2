module ff_e_c_rn(
    input D,
    input E,
    input CP,
    input CDN,
    output Q
);
endmodule
