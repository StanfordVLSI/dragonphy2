module termination (
	input VinP,
	input VinN,
	input Vcm
);
endmodule