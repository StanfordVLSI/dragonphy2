package test_pack;

	localparam real full_rate = 16e9;

endpackage
