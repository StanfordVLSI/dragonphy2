module ff_c_rn(
    input D,
    input CP,
    input CDN,
    output Q
);
endmodule
