
module inv_v2t_4_fixed (input in, output out );
assign out = ~(in);
endmodule

