module inv_xc (
    input in,
    output out
);
endmodule

