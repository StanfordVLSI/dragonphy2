module input_buffer_inv (
    input inp,
    input inm,
    input pd,
    output clk,
    output clk_b
);
endmodule