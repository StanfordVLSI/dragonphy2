
module dcdl_coarse ( out, in, thm );
  input [30:0] thm;
  input in;
  output out;
  wire   dr0, dm0;
  wire   [30:0] dm;
  wire   [29:0] dr;
  wire   [30:0] df;
  wire   [30:0] thm_b;

  n_and I89_0_ ( .in1(dr[0]), .in2(dm[0]), .out(dr0) );
  n_and I89_1_ ( .in1(dr[1]), .in2(dm[1]), .out(dr[0]) );
  n_and I89_2_ ( .in1(dr[2]), .in2(dm[2]), .out(dr[1]) );
  n_and I89_3_ ( .in1(dr[3]), .in2(dm[3]), .out(dr[2]) );
  n_and I89_4_ ( .in1(dr[4]), .in2(dm[4]), .out(dr[3]) );
  n_and I89_5_ ( .in1(dr[5]), .in2(dm[5]), .out(dr[4]) );
  n_and I89_6_ ( .in1(dr[6]), .in2(dm[6]), .out(dr[5]) );
  n_and I89_7_ ( .in1(dr[7]), .in2(dm[7]), .out(dr[6]) );
  n_and I89_8_ ( .in1(dr[8]), .in2(dm[8]), .out(dr[7]) );
  n_and I89_9_ ( .in1(dr[9]), .in2(dm[9]), .out(dr[8]) );
  n_and I89_10_ ( .in1(dr[10]), .in2(dm[10]), .out(dr[9]) );
  n_and I89_11_ ( .in1(dr[11]), .in2(dm[11]), .out(dr[10]) );
  n_and I89_12_ ( .in1(dr[12]), .in2(dm[12]), .out(dr[11]) );
  n_and I89_13_ ( .in1(dr[13]), .in2(dm[13]), .out(dr[12]) );
  n_and I89_14_ ( .in1(dr[14]), .in2(dm[14]), .out(dr[13]) );
  n_and I89_15_ ( .in1(dr[15]), .in2(dm[15]), .out(dr[14]) );
  n_and I89_16_ ( .in1(dr[16]), .in2(dm[16]), .out(dr[15]) );
  n_and I89_17_ ( .in1(dr[17]), .in2(dm[17]), .out(dr[16]) );
  n_and I89_18_ ( .in1(dr[18]), .in2(dm[18]), .out(dr[17]) );
  n_and I89_19_ ( .in1(dr[19]), .in2(dm[19]), .out(dr[18]) );
  n_and I89_20_ ( .in1(dr[20]), .in2(dm[20]), .out(dr[19]) );
  n_and I89_21_ ( .in1(dr[21]), .in2(dm[21]), .out(dr[20]) );
  n_and I89_22_ ( .in1(dr[22]), .in2(dm[22]), .out(dr[21]) );
  n_and I89_23_ ( .in1(dr[23]), .in2(dm[23]), .out(dr[22]) );
  n_and I89_24_ ( .in1(dr[24]), .in2(dm[24]), .out(dr[23]) );
  n_and I89_25_ ( .in1(dr[25]), .in2(dm[25]), .out(dr[24]) );
  n_and I89_26_ ( .in1(dr[26]), .in2(dm[26]), .out(dr[25]) );
  n_and I89_27_ ( .in1(dr[27]), .in2(dm[27]), .out(dr[26]) );
  n_and I89_28_ ( .in1(dr[28]), .in2(dm[28]), .out(dr[27]) );
  n_and I89_29_ ( .in1(dr[29]), .in2(dm[29]), .out(dr[28]) );
  n_and I89_30_ ( .in1(1'b1), .in2(dm[30]), .out(dr[29]) );
  n_and I88_0_ ( .in1(thm_b[1]), .in2(df[0]), .out(dm[0]) );
  n_and I88_1_ ( .in1(thm_b[2]), .in2(df[1]), .out(dm[1]) );
  n_and I88_2_ ( .in1(thm_b[3]), .in2(df[2]), .out(dm[2]) );
  n_and I88_3_ ( .in1(thm_b[4]), .in2(df[3]), .out(dm[3]) );
  n_and I88_4_ ( .in1(thm_b[5]), .in2(df[4]), .out(dm[4]) );
  n_and I88_5_ ( .in1(thm_b[6]), .in2(df[5]), .out(dm[5]) );
  n_and I88_6_ ( .in1(thm_b[7]), .in2(df[6]), .out(dm[6]) );
  n_and I88_7_ ( .in1(thm_b[8]), .in2(df[7]), .out(dm[7]) );
  n_and I88_8_ ( .in1(thm_b[9]), .in2(df[8]), .out(dm[8]) );
  n_and I88_9_ ( .in1(thm_b[10]), .in2(df[9]), .out(dm[9]) );
  n_and I88_10_ ( .in1(thm_b[11]), .in2(df[10]), .out(dm[10]) );
  n_and I88_11_ ( .in1(thm_b[12]), .in2(df[11]), .out(dm[11]) );
  n_and I88_12_ ( .in1(thm_b[13]), .in2(df[12]), .out(dm[12]) );
  n_and I88_13_ ( .in1(thm_b[14]), .in2(df[13]), .out(dm[13]) );
  n_and I88_14_ ( .in1(thm_b[15]), .in2(df[14]), .out(dm[14]) );
  n_and I88_15_ ( .in1(thm_b[16]), .in2(df[15]), .out(dm[15]) );
  n_and I88_16_ ( .in1(thm_b[17]), .in2(df[16]), .out(dm[16]) );
  n_and I88_17_ ( .in1(thm_b[18]), .in2(df[17]), .out(dm[17]) );
  n_and I88_18_ ( .in1(thm_b[19]), .in2(df[18]), .out(dm[18]) );
  n_and I88_19_ ( .in1(thm_b[20]), .in2(df[19]), .out(dm[19]) );
  n_and I88_20_ ( .in1(thm_b[21]), .in2(df[20]), .out(dm[20]) );
  n_and I88_21_ ( .in1(thm_b[22]), .in2(df[21]), .out(dm[21]) );
  n_and I88_22_ ( .in1(thm_b[23]), .in2(df[22]), .out(dm[22]) );
  n_and I88_23_ ( .in1(thm_b[24]), .in2(df[23]), .out(dm[23]) );
  n_and I88_24_ ( .in1(thm_b[25]), .in2(df[24]), .out(dm[24]) );
  n_and I88_25_ ( .in1(thm_b[26]), .in2(df[25]), .out(dm[25]) );
  n_and I88_26_ ( .in1(thm_b[27]), .in2(df[26]), .out(dm[26]) );
  n_and I88_27_ ( .in1(thm_b[28]), .in2(df[27]), .out(dm[27]) );
  n_and I88_28_ ( .in1(thm_b[29]), .in2(df[28]), .out(dm[28]) );
  n_and I88_29_ ( .in1(thm_b[30]), .in2(df[29]), .out(dm[29]) );
  n_and I88_30_ ( .in1(1'b1), .in2(df[30]), .out(dm[30]) );
  n_and I85 ( .in1(thm_b[0]), .in2(in), .out(dm0) );
  n_and I87_0_ ( .in1(thm[0]), .in2(in), .out(df[0]) );
  n_and I87_1_ ( .in1(thm[1]), .in2(df[0]), .out(df[1]) );
  n_and I87_2_ ( .in1(thm[2]), .in2(df[1]), .out(df[2]) );
  n_and I87_3_ ( .in1(thm[3]), .in2(df[2]), .out(df[3]) );
  n_and I87_4_ ( .in1(thm[4]), .in2(df[3]), .out(df[4]) );
  n_and I87_5_ ( .in1(thm[5]), .in2(df[4]), .out(df[5]) );
  n_and I87_6_ ( .in1(thm[6]), .in2(df[5]), .out(df[6]) );
  n_and I87_7_ ( .in1(thm[7]), .in2(df[6]), .out(df[7]) );
  n_and I87_8_ ( .in1(thm[8]), .in2(df[7]), .out(df[8]) );
  n_and I87_9_ ( .in1(thm[9]), .in2(df[8]), .out(df[9]) );
  n_and I87_10_ ( .in1(thm[10]), .in2(df[9]), .out(df[10]) );
  n_and I87_11_ ( .in1(thm[11]), .in2(df[10]), .out(df[11]) );
  n_and I87_12_ ( .in1(thm[12]), .in2(df[11]), .out(df[12]) );
  n_and I87_13_ ( .in1(thm[13]), .in2(df[12]), .out(df[13]) );
  n_and I87_14_ ( .in1(thm[14]), .in2(df[13]), .out(df[14]) );
  n_and I87_15_ ( .in1(thm[15]), .in2(df[14]), .out(df[15]) );
  n_and I87_16_ ( .in1(thm[16]), .in2(df[15]), .out(df[16]) );
  n_and I87_17_ ( .in1(thm[17]), .in2(df[16]), .out(df[17]) );
  n_and I87_18_ ( .in1(thm[18]), .in2(df[17]), .out(df[18]) );
  n_and I87_19_ ( .in1(thm[19]), .in2(df[18]), .out(df[19]) );
  n_and I87_20_ ( .in1(thm[20]), .in2(df[19]), .out(df[20]) );
  n_and I87_21_ ( .in1(thm[21]), .in2(df[20]), .out(df[21]) );
  n_and I87_22_ ( .in1(thm[22]), .in2(df[21]), .out(df[22]) );
  n_and I87_23_ ( .in1(thm[23]), .in2(df[22]), .out(df[23]) );
  n_and I87_24_ ( .in1(thm[24]), .in2(df[23]), .out(df[24]) );
  n_and I87_25_ ( .in1(thm[25]), .in2(df[24]), .out(df[25]) );
  n_and I87_26_ ( .in1(thm[26]), .in2(df[25]), .out(df[26]) );
  n_and I87_27_ ( .in1(thm[27]), .in2(df[26]), .out(df[27]) );
  n_and I87_28_ ( .in1(thm[28]), .in2(df[27]), .out(df[28]) );
  n_and I87_29_ ( .in1(thm[29]), .in2(df[28]), .out(df[29]) );
  n_and I87_30_ ( .in1(thm[30]), .in2(df[29]), .out(df[30]) );
  n_and I84 ( .in1(dr0), .in2(dm0), .out(out) );
  inv I83_0_ ( .in(thm[0]), .out(thm_b[0]) );
  inv I83_1_ ( .in(thm[1]), .out(thm_b[1]) );
  inv I83_2_ ( .in(thm[2]), .out(thm_b[2]) );
  inv I83_3_ ( .in(thm[3]), .out(thm_b[3]) );
  inv I83_4_ ( .in(thm[4]), .out(thm_b[4]) );
  inv I83_5_ ( .in(thm[5]), .out(thm_b[5]) );
  inv I83_6_ ( .in(thm[6]), .out(thm_b[6]) );
  inv I83_7_ ( .in(thm[7]), .out(thm_b[7]) );
  inv I83_8_ ( .in(thm[8]), .out(thm_b[8]) );
  inv I83_9_ ( .in(thm[9]), .out(thm_b[9]) );
  inv I83_10_ ( .in(thm[10]), .out(thm_b[10]) );
  inv I83_11_ ( .in(thm[11]), .out(thm_b[11]) );
  inv I83_12_ ( .in(thm[12]), .out(thm_b[12]) );
  inv I83_13_ ( .in(thm[13]), .out(thm_b[13]) );
  inv I83_14_ ( .in(thm[14]), .out(thm_b[14]) );
  inv I83_15_ ( .in(thm[15]), .out(thm_b[15]) );
  inv I83_16_ ( .in(thm[16]), .out(thm_b[16]) );
  inv I83_17_ ( .in(thm[17]), .out(thm_b[17]) );
  inv I83_18_ ( .in(thm[18]), .out(thm_b[18]) );
  inv I83_19_ ( .in(thm[19]), .out(thm_b[19]) );
  inv I83_20_ ( .in(thm[20]), .out(thm_b[20]) );
  inv I83_21_ ( .in(thm[21]), .out(thm_b[21]) );
  inv I83_22_ ( .in(thm[22]), .out(thm_b[22]) );
  inv I83_23_ ( .in(thm[23]), .out(thm_b[23]) );
  inv I83_24_ ( .in(thm[24]), .out(thm_b[24]) );
  inv I83_25_ ( .in(thm[25]), .out(thm_b[25]) );
  inv I83_26_ ( .in(thm[26]), .out(thm_b[26]) );
  inv I83_27_ ( .in(thm[27]), .out(thm_b[27]) );
  inv I83_28_ ( .in(thm[28]), .out(thm_b[28]) );
  inv I83_29_ ( .in(thm[29]), .out(thm_b[29]) );
  inv I83_30_ ( .in(thm[30]), .out(thm_b[30]) );
endmodule

