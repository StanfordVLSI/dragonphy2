module tm_stall ();
endmodule
