
module inv_arb_fixed (input in, output out );
assign out = ~(in);
endmodule

