
module inv_v2t_1_fixed (input in, output out );
assign out = ~(in);
endmodule

