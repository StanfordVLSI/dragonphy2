module input_buffer (
	input inp,
	input inn,
	input en,
	input in_aux,
	input sel_in,
	input bypass_div,
	input [2:0] ndiv,
	input en_meas,

	output out,
	output out_meas
);
endmodule