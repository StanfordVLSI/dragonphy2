
module CS_cell (input Vbias, input CTRL, input CS_DRN);
endmodule


