module vio (
    output wire logic emu_rst,
    output wire logic rst_user,
    input wire logic [63:0] number,
    input wire logic clk
);

endmodule
