
module inv_bld_2_fixed (input in, output out );
assign out = ~(in);
endmodule

