`define ANALOG_INPUT inout wire
`define ANALOG_OUTPUT inout wire

`define DECL_ANALOG(x) wire x;
