module inv_skewed (
    input in,
    output out
);
endmodule

