module ff_cn_sn_rn(
    input D,
    input CPN,
    input CDN,
    input SDN,
    output Q
);
endmodule
