module TS1N16FFCLLSBLVTC1024X144M4SW (
	input CLK,
	input CEB,
	input WEB,
	input [9:0] A,
	input [143:0] D,
	output [143:0] Q,
	input [143:0] BWEB,
	input [1:0] RTSEL,
	input [1:0] WTSEL
);
endmodule