module sram_144_1024_freepdk45 (
	input clk0,
	input csb0,
	input web0,
	input [9:0] addr0,
	input [143:0] din0,
	output [143:0] dout0
);
endmodule
