
module inv_v2t_0_fixed (input in, output out );
assign out = ~(in);
endmodule

