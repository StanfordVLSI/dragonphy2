module tri_buff (
    input in,
    input en,
    output out
);

bufif1(out,in,en);

endmodule




