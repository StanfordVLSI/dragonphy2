module ff_e_c_rn(
    input D,
    input E,
    input CP,
    output Q,
    input CDN,
);
endmodule
