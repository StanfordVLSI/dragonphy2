module BUFG (
    output wire logic O,
    input wire logic I
);

    assign O = I;

endmodule
