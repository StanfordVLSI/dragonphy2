
module inv (input in, output out );
assign out = ~(in);
endmodule

