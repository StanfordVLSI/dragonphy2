
module inv_0_fixed (input in, output out );
assign out = ~(in);
endmodule

