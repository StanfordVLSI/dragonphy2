module inv_3 (
    input in,
    output out
);
endmodule

