
module inv_1_fixed (input in, output out );
assign out = ~(in);
endmodule

