`include "mLingua_pwl.vh"

`default_nettype none

module termination import const_pack::* ; #(
) (
	input pwl VinP,
	input pwl VinN,
	input real Vcm
);

endmodule

`default_nettype wire