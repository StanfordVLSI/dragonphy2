module ff_c_sn_rn(
    input D,
    input CP,
    output Q,
    input CDN,
);
endmodule
