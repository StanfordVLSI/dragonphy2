
module inv_PI_2_fixed (input in, output out );
assign out = ~(in);
endmodule

