
module inv_v2t_3_fixed (input in, output out );
assign out = ~(in);
endmodule

