
module inv_bld_1_fixed (input in, output out );
assign out = ~(in);
endmodule

