module inv_4 (
    input in,
    output out
);
endmodule

