module mmcm (
    input wire logic ext_clk,
    output var logic emu_clk_2x
);

    // instantiate clock wizard here...

endmodule

