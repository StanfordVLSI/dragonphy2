module test;
	initial begin
		$display("Hello world!");
		$finish;
	end
endmodule
