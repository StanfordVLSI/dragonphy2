
module inv_PI_1_fixed (input in, output out );
assign out = ~(in);
endmodule

