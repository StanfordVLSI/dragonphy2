
module inv_PI (input in, output out );
assign out = ~(in);
endmodule

