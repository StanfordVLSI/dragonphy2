module ff_cn_sn_rn(
    input D,
    input CPN,
    output Q,
    input CDN,
    input SDN
);
endmodule
