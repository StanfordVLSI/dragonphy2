
module inv_5_fixed (input in, output out );
assign out = ~(in);
endmodule

