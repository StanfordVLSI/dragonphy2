interface analog_if ();
    real value;
endinterface

`define ANALOG_INPUT interface
`define ANALOG_OUTPUT interface

`define DECL_ANALOG(x) analog_if x ()
