module termination (
	input pwl VinP,
	input pwl VinN,
	input real Vcm
);
endmodule