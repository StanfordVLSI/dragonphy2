module inc_delay (
    input in,
    input inc_del,
    output out
);
endmodule