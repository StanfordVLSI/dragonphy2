module ff(
    input D,
    input CPN,
    output Q,
    input CDN,
    input SDN
);
endmodule
