module input_buffer (
	input inp,
	input inm,
	input pd,
	output clk,
	output clk_b
);

    assign clk = 1'b0;
    assign clk_b = 1'b0;

endmodule
